-- =====================================================
-- 📦 Package com tipo personalizado
-- =====================================================
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package Types is
    type array_3X7bits is array (0 to 6) of std_logic_vector(2 downto 0);
end package Types;

package body Types is
end package body Types;
